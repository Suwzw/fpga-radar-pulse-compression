//-----------------------------------------------------------------------------
// Module: clt_noise_generator
//
// Description:
//   使用中央极限定理生成近似高斯白噪声。
//   它例化N个LFSR，并将它们的单比特输出相加。
//-----------------------------------------------------------------------------
module clt_noise_generator #(
    parameter NUM_LFSRS = 12 // 使用的LFSR数量
) (
    input  wire clk,
    input  wire rst_n,

    // 输出的噪声样本，是有符号数
    // 范围是 [-6, +6] (对于NUM_LFSRS=12)
    output wire signed [4:0] noise_out
);

    // 用于连接所有LFSR输出比特的线网
    wire [NUM_LFSRS-1:0] lfsr_bits;

    // 使用Verilog的generate语句，批量例化12个LFSR
    // 这是非常强大和可扩展的写法
    genvar i;
    generate
        for (i = 0; i < NUM_LFSRS; i = i + 1) begin : lfsr_inst
            // 关键：为每个LFSR提供一个不同的、非零的初始种子
            // 这里我们简单地使用一个递增的值
            lfsr #(
                .WIDTH(16),
                .INITIAL_SEED(16'h1234 + i) 
            ) u_lfsr (
                .clk(clk),
                .rst_n(rst_n),
                .random_bit_out(lfsr_bits[i])
            );
        end
    endgenerate

    //--- 求和与均值调整 ---

    // 1. 求和
    // 对12个比特(0或1)求和，结果范围是[0, 12]
    // 需要 ceil(log2(12+1)) = 4 位来表示这个和
    wire [3:0] sum_unsigned;
    
    // 用一个assign语句实现并行加法器树
    assign sum_unsigned = lfsr_bits[0]  + lfsr_bits[1]  + lfsr_bits[2]  + lfsr_bits[3] +
                        lfsr_bits[4]  + lfsr_bits[5]  + lfsr_bits[6]  + lfsr_bits[7] +
                        lfsr_bits[8]  + lfsr_bits[9]  + lfsr_bits[10] + lfsr_bits[11];
    
    // 2. 均值调整 (减去均值，使其变为零均值噪声)
    // 12个LFSR输出的和的期望值(均值)是 12 * 0.5 = 6
    // 我们将和减去6，使得新序列的均值为0。
    // 原始和范围: [0, 1, ..., 12]
    // 减6后范围: [-6, -5, ..., 6]
    // 这个范围需要5位有符号数来表示
    localparam MEAN_ADJUST = NUM_LFSRS / 2;
    
    assign noise_out = sum_unsigned - MEAN_ADJUST;

endmodule