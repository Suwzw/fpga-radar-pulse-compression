`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: Interpolate
// Description: R����ֵģ�顣���յ�һ��������Ч����ʱ�����R�������㣬
//              ��һ��Ϊ�������ݱ�������R-1��Ϊ�㡣
//              �ȴ���һ����ʱ���ڿ���״̬��
//////////////////////////////////////////////////////////////////////////////////
module Interpolate #(
    parameter R = 4,               // ��ֵ������Ĭ��4����ֵ
    parameter INPUT_WIDTH = 14,    // ��������λ��
    parameter OUTPUT_WIDTH = 22    // �������λ��
)(
    input                       rst,        // ��λ�źţ��ߵ�ƽ��Ч
    input                       clk,        // ʱ���ź�
    input  signed [INPUT_WIDTH-1:0] Xin,    // ������������
    input                       Xin_valid,  // ����������Ч�ź�
    output reg signed [OUTPUT_WIDTH-1:0] Xout,  // �����������
    output reg                  Xout_valid  // ���������Ч�ź�
);

    reg [31:0] count = 0;
    reg busy = 0;                   // ��ǵ�ǰ�Ƿ��������ֵ����
    reg signed [OUTPUT_WIDTH-1:0] sample_buffer;

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            count <= 0;
            busy <= 0;
            Xout <= 0;
            Xout_valid <= 0;
            sample_buffer <= 0;
        end else begin
            Xout_valid <= 0; // Ĭ�ϱ������������Ч��������������
            if (busy) begin
                // �����æ�������ֵ����
                if (count < R) begin
                    // �����count������
                    if (count == 0) begin
                        // ��һ���������Ϊ�洢���������㣬������չ��OUTPUT_WIDTH
                        Xout <= {{(OUTPUT_WIDTH-INPUT_WIDTH){sample_buffer[INPUT_WIDTH-1]}}, sample_buffer[INPUT_WIDTH-1:0]};
                    end else begin
                        // ʣ���R-1�����Ϊ0
                        Xout <= 0;
                    end
                    Xout_valid <= 1;
                    count <= count + 1;
                end else begin
                    // �������R���㣬������еȴ���һ����������
                    busy <= 0;
                end
            end else begin
                // ����״̬�µȴ��µ�������Ч����
                if (Xin_valid) begin
                    // �洢�������㣬׼�����R����
                    sample_buffer <= {{(OUTPUT_WIDTH-INPUT_WIDTH){Xin[INPUT_WIDTH-1]}}, Xin};
                    count <= 0;
                    busy <= 1;
                end
            end
        end
    end
endmodule
