`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Module Name: Decimate
// Description: R����ȡģ�飬ͨ������R���Ƴ�ȡ����
//////////////////////////////////////////////////////////////////////////////////

module Decimate #(
    parameter R = 5,               // ��ȡ�����������ɸ�����Ҫ����
    parameter DATA_WIDTH = 22      // �����������λ���ɸ���ʵ���������
)(
    input               rst,       // ��λ�źţ��ߵ�ƽ��Ч
    input               clk,       // FPGAϵͳʱ��
    input  signed [DATA_WIDTH-1:0] Iin,  // ��������
    output signed [DATA_WIDTH-1:0] dout, // �������(��ȡ��)
    output              rdy        // ������Ч����ź�
);

    // ���������ڿ��ƺ�ʱ�������
    // ����������0������R-1ʱ������ݣ�Ȼ������
    reg [$clog2(R)-1:0] c = 0;      // ���������ȡ����R�Ĵ�С
    reg signed [DATA_WIDTH-1:0] dout_tem = 0; // �������
    reg rdy_tem = 0;                 // ������Ч�ź�

    // ��λ�߼�����ʼ�����мĴ���
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            // �����λ�ź�Ϊ�ߣ����мĴ�������
            c <= 0;
            dout_tem <= {DATA_WIDTH{1'b0}}; // ��λʱ��������
            rdy_tem <= 1'b0;                // ������Ч�ź�����
        end else begin
            // �Ǹ�λ״̬��ִ�г�ȡ�߼�
            if (c == R-1) begin
                // �����ﵽR-1ʱ�����������Ч
                rdy_tem <= 1'b1;
                dout_tem <= Iin;  // �洢�������ݵ�������ݼĴ���
                c <= 0;            // ���ü�����
            end else begin
                // ������δ�ﵽR-1ʱ�����������
                rdy_tem <= 1'b0;
                c <= c + 1;        // ��������1
            end
        end
    end

    // ��������������Ľ����������ź�
    assign dout = dout_tem; // �����ȡ�������
    assign rdy  = rdy_tem;  // ���������Ч�ź�

endmodule
