`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: MultCIC (Corrected Control Signal Version)
// Description: CIC�˲�������ģ�飬��������ֵģʽ�µĿ����ź�bug
//////////////////////////////////////////////////////////////////////////////////
module MultCIC #(
    parameter MODE = "DEC",      // "DEC" �� "INT" ģʽ��ѡ����ģʽ
    parameter R = 5,             // ��ȡ���ֵ�ı�����Ӱ�������
    parameter D = 3,             // ���ּ���������CIC�˲����ļ���
    parameter INPUT_WIDTH = 14,  // ��������λ��
    parameter OUTPUT_WIDTH = 22  // �������λ��
)(
    input        rst,            // ��λ�źţ��ߵ�ƽ��Ч
    input        clk,            // ʱ���ź�
    input  [INPUT_WIDTH-1:0] Xin, // ��������
    // --- START: �����޸� ---
    input        Xin_valid,      // Ϊ��ֵģʽ������������Ч�ź�
    // --- END: �����޸� ---
    output [OUTPUT_WIDTH-1:0] Yout, // �������
    output        rdy            // ������Чָʾ�ź�
);


    // �м��ź�
    wire signed [OUTPUT_WIDTH-1:0] Intout;   // ����ģ���������
    wire signed [OUTPUT_WIDTH-1:0] dout;     // ��ȡģ���������
    wire ND;  // ������Ч�ź�


    // ���ɲ�ͬģʽ�µ�ģ��ʵ��
    generate
        // ���ѡ���ȡģʽ��"DEC"������ִ�����´���
        if (MODE == "DEC") begin : DEC_MODE

            // 1. ʵ����������ģ��
            Integrated #(
                .D(D),                // ���ּ���
                .INPUT_WIDTH(INPUT_WIDTH),  // ��������λ��
                .OUTPUT_WIDTH(OUTPUT_WIDTH) // �������λ��
            ) U_Int (
                .rst(rst),            // ��λ�ź�
                .clk(clk),            // ʱ���ź�
                .Xin(Xin),            // ��������
                .Intout(Intout)       // �����������
            );



            // 2. ʵ������ȡģ��
            // ��ȡģ�����Rֵ������ȡ�ı�������С������ݵ�����
            Decimate #(
                .R(R),                // ��ȡ����
                .DATA_WIDTH(OUTPUT_WIDTH)  // ������ݿ��
            ) U_Dec (
                .rst(rst),            // ��λ�ź�
                .clk(clk),            // ʱ���ź�
                .Iin(Intout),         // ��������
                .dout(dout),          // ��ȡ�������
                .rdy(ND)              // ������Чָʾ�ź�
            );



            // 3. ʵ������״�˲�����Comb�������в�ֲ���
            Comb #(
                .D(D),                        // ��ּ���
                .DATA_WIDTH(OUTPUT_WIDTH)     // ������ݿ��
            ) U_Comb (
                .rst(rst),                    // ��λ�ź�
                .clk(clk),                    // ʱ���ź�
                .ND(ND),                      // ������Ч�ź�
                .Xin(dout),                   // ��������
                .Yout(Yout)                   // ��״�˲������������
            );

            // ���������Ч�ź�
            assign rdy = ND;

        end else if (MODE == "INT") begin : INT_MODE

            // 1. ��ֵģʽ�µ���״�˲�����Comb��
            wire signed [OUTPUT_WIDTH-1:0] comb_out;    // ��״�˲����������
            wire signed [OUTPUT_WIDTH-1:0] interp_out;  // ��ֵ�������
            wire interp_rdy;                           // ��ֵģ���������Ч�ź�


            // --- START: �����޸� ---
            // ��״�˲���ֻ��������Чʱ��ʹ��
            Comb #(
                .D(D),                        // ��ּ���
                .DATA_WIDTH(OUTPUT_WIDTH)     // ������ݿ��
            ) U_Comb_int (
                .rst(rst),                    // ��λ�ź�
                .clk(clk),                    // ʱ���ź�
                .ND(Xin_valid),               // <<--- �޸ĵ㣺ʹ���ⲿ��Ч�ź�
                .Xin({{(OUTPUT_WIDTH-INPUT_WIDTH){Xin[INPUT_WIDTH-1]}}, Xin}),  // �����źŷ�����չ
                .Yout(comb_out)               // ��״�˲��������
            );


            // 2. ʵ������ֵģ�飨Interpolate��
            // ���ݲ�ֵ����R��������в���R-1�����
            Interpolate #(
                .R(R),                // ��ֵ����
                .INPUT_WIDTH(OUTPUT_WIDTH),  // ��������λ��
                .OUTPUT_WIDTH(OUTPUT_WIDTH)  // �������λ��
            ) U_Interp (
                .rst(rst),            // ��λ�ź�
                .clk(clk),            // ʱ���ź�
                .Xin(comb_out),       // ���ݸ���ֵģ�������
                .Xin_valid(Xin_valid), // <<--- �޸ĵ㣺ʹ���ⲿ��Ч�ź�
                .Xout(interp_out),    // ��ֵ�������
                .Xout_valid(interp_rdy) // ��ֵ��Ч�ź�
            );
            // --- END: �����޸� ---
            

            // 3. ��ֵ�����ݽ��������
            Integrated #(
                .D(D),                // ���ּ���
                .INPUT_WIDTH(OUTPUT_WIDTH),  // ��������λ��
                .OUTPUT_WIDTH(OUTPUT_WIDTH) // �������λ��
            ) U_Int_int (
                .rst(rst),            // ��λ�ź�
                .clk(clk),            // ʱ���ź�
                .Xin(interp_out[OUTPUT_WIDTH-1:0]),  // ��ֵ������ݣ�������Ҫ�ضϣ�
                .Intout(Yout)         // �������������
            );

            // �����ֵ������Ч�ź�
            assign rdy = interp_rdy;

        end else begin : DEFAULT_MODE
            // Ĭ��ģʽ����MODE�Ȳ���"DEC"Ҳ����"INT"ʱ�������Ч
            assign Yout = {OUTPUT_WIDTH{1'b0}}; // ���ȫ0
            assign rdy = 1'b0; // �����Ч�ź�
        end
    endgenerate

endmodule
